module SR(
);

  // TODO

endmodule